module MeshWrapper
(
    input clk,
    input rst,

    input [16-1:0] in_input_0_payload_discriminant,
    input [128-1:0] in_input_0_payload_Some_0_a_0,
    input [16-1:0] in_input_1_0_payload_discriminant,
    input [320-1:0] in_input_1_0_payload_Some_0_b_0,
    input [320-1:0] in_input_1_0_payload_Some_0_d_0,
    input [16-1:0] in_input_1_1_payload_discriminant,
    input [48-1:0] in_input_1_1_payload_Some_0_id,
    input [16-1:0] in_input_1_1_payload_Some_0_last,
    input [16-1:0] in_input_1_1_payload_Some_0_control_dataflow_discriminant,
    input [16-1:0] in_input_1_1_payload_Some_0_control_propagate_discriminant,
    input [80-1:0] in_input_1_1_payload_Some_0_control_shift,
    input [16-1:0] in_input_1_1_payload_Some_0_bad_dataflow,

    output [16-1:0] out_output_0_payload_discriminant, // DontCare
    output [128-1:0] out_output_0_payload_Some_0_a_0,    // DontCare
    output [16-1:0] out_output_1_0_payload_discriminant,
    output [320-1:0] out_output_1_0_payload_Some_0_b_0,
    output [320-1:0] out_output_1_0_payload_Some_0_d_0,
    output [16-1:0] out_output_1_1_payload_discriminant,
    output [48-1:0] out_output_1_1_payload_Some_0_id,
    output [16-1:0] out_output_1_1_payload_Some_0_last,
    output [16-1:0] out_output_1_1_payload_Some_0_control_dataflow_discriminant,
    output [16-1:0] out_output_1_1_payload_Some_0_control_propagate_discriminant, // DontCare
    output [80-1:0] out_output_1_1_payload_Some_0_control_shift, // DontCare
    output [16-1:0] out_output_1_1_payload_Some_0_bad_dataflow   // DontCare
);
    wire io_out_valid_0_0;
    wire io_out_control_0_0_dataflow;
    wire [2:0] io_out_id_0_0;
    wire io_out_last_0_0;

    Mesh mesh_inst(
        .clock(clk),
        .reset(rst),

        .io_in_a_0_0(in_input_0_payload_Some_0_a_0[0*8 +: 8]),
        .io_in_a_1_0(in_input_0_payload_Some_0_a_0[1*8 +: 8]),
        .io_in_a_2_0(in_input_0_payload_Some_0_a_0[2*8 +: 8]),
        .io_in_a_3_0(in_input_0_payload_Some_0_a_0[3*8 +: 8]),
        .io_in_a_4_0(in_input_0_payload_Some_0_a_0[4*8 +: 8]),
        .io_in_a_5_0(in_input_0_payload_Some_0_a_0[5*8 +: 8]),
        .io_in_a_6_0(in_input_0_payload_Some_0_a_0[6*8 +: 8]),
        .io_in_a_7_0(in_input_0_payload_Some_0_a_0[7*8 +: 8]),
        .io_in_a_8_0(in_input_0_payload_Some_0_a_0[8*8 +: 8]),
        .io_in_a_9_0(in_input_0_payload_Some_0_a_0[9*8 +: 8]),
        .io_in_a_10_0(in_input_0_payload_Some_0_a_0[10*8 +: 8]),
        .io_in_a_11_0(in_input_0_payload_Some_0_a_0[11*8 +: 8]),
        .io_in_a_12_0(in_input_0_payload_Some_0_a_0[12*8 +: 8]),
        .io_in_a_13_0(in_input_0_payload_Some_0_a_0[13*8 +: 8]),
        .io_in_a_14_0(in_input_0_payload_Some_0_a_0[14*8 +: 8]),
        .io_in_a_15_0(in_input_0_payload_Some_0_a_0[15*8 +: 8]),

        .io_in_b_0_0(in_input_1_0_payload_Some_0_b_0[0*20 +: 20]),
        .io_in_b_1_0(in_input_1_0_payload_Some_0_b_0[1*20 +: 20]),
        .io_in_b_2_0(in_input_1_0_payload_Some_0_b_0[2*20 +: 20]),
        .io_in_b_3_0(in_input_1_0_payload_Some_0_b_0[3*20 +: 20]),
        .io_in_b_4_0(in_input_1_0_payload_Some_0_b_0[4*20 +: 20]),
        .io_in_b_5_0(in_input_1_0_payload_Some_0_b_0[5*20 +: 20]),
        .io_in_b_6_0(in_input_1_0_payload_Some_0_b_0[6*20 +: 20]),
        .io_in_b_7_0(in_input_1_0_payload_Some_0_b_0[7*20 +: 20]),
        .io_in_b_8_0(in_input_1_0_payload_Some_0_b_0[8*20 +: 20]),
        .io_in_b_9_0(in_input_1_0_payload_Some_0_b_0[9*20 +: 20]),
        .io_in_b_10_0(in_input_1_0_payload_Some_0_b_0[10*20 +: 20]),
        .io_in_b_11_0(in_input_1_0_payload_Some_0_b_0[11*20 +: 20]),
        .io_in_b_12_0(in_input_1_0_payload_Some_0_b_0[12*20 +: 20]),
        .io_in_b_13_0(in_input_1_0_payload_Some_0_b_0[13*20 +: 20]),
        .io_in_b_14_0(in_input_1_0_payload_Some_0_b_0[14*20 +: 20]),
        .io_in_b_15_0(in_input_1_0_payload_Some_0_b_0[15*20 +: 20]),

        .io_in_d_0_0(in_input_1_0_payload_Some_0_d_0[0*20 +: 20]),
        .io_in_d_1_0(in_input_1_0_payload_Some_0_d_0[1*20 +: 20]),
        .io_in_d_2_0(in_input_1_0_payload_Some_0_d_0[2*20 +: 20]),
        .io_in_d_3_0(in_input_1_0_payload_Some_0_d_0[3*20 +: 20]),
        .io_in_d_4_0(in_input_1_0_payload_Some_0_d_0[4*20 +: 20]),
        .io_in_d_5_0(in_input_1_0_payload_Some_0_d_0[5*20 +: 20]),
        .io_in_d_6_0(in_input_1_0_payload_Some_0_d_0[6*20 +: 20]),
        .io_in_d_7_0(in_input_1_0_payload_Some_0_d_0[7*20 +: 20]),
        .io_in_d_8_0(in_input_1_0_payload_Some_0_d_0[8*20 +: 20]),
        .io_in_d_9_0(in_input_1_0_payload_Some_0_d_0[9*20 +: 20]),
        .io_in_d_10_0(in_input_1_0_payload_Some_0_d_0[10*20 +: 20]),
        .io_in_d_11_0(in_input_1_0_payload_Some_0_d_0[11*20 +: 20]),
        .io_in_d_12_0(in_input_1_0_payload_Some_0_d_0[12*20 +: 20]),
        .io_in_d_13_0(in_input_1_0_payload_Some_0_d_0[13*20 +: 20]),
        .io_in_d_14_0(in_input_1_0_payload_Some_0_d_0[14*20 +: 20]),
        .io_in_d_15_0(in_input_1_0_payload_Some_0_d_0[15*20 +: 20]),

        .io_in_control_0_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[0]),
        .io_in_control_0_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[0]),
        .io_in_control_0_0_shift(in_input_1_1_payload_Some_0_control_shift[0*5 +: 5]),
        .io_in_control_1_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[1]),
        .io_in_control_1_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[1]),
        .io_in_control_1_0_shift(in_input_1_1_payload_Some_0_control_shift[1*5 +: 5]),
        .io_in_control_2_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[2]),
        .io_in_control_2_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[2]),
        .io_in_control_2_0_shift(in_input_1_1_payload_Some_0_control_shift[2*5 +: 5]),
        .io_in_control_3_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[3]),
        .io_in_control_3_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[3]),
        .io_in_control_3_0_shift(in_input_1_1_payload_Some_0_control_shift[3*5 +: 5]),
        .io_in_control_4_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[4]),
        .io_in_control_4_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[4]),
        .io_in_control_4_0_shift(in_input_1_1_payload_Some_0_control_shift[4*5 +: 5]),
        .io_in_control_5_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[5]),
        .io_in_control_5_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[5]),
        .io_in_control_5_0_shift(in_input_1_1_payload_Some_0_control_shift[5*5 +: 5]),
        .io_in_control_6_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[6]),
        .io_in_control_6_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[6]),
        .io_in_control_6_0_shift(in_input_1_1_payload_Some_0_control_shift[6*5 +: 5]),
        .io_in_control_7_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[7]),
        .io_in_control_7_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[7]),
        .io_in_control_7_0_shift(in_input_1_1_payload_Some_0_control_shift[7*5 +: 5]),
        .io_in_control_8_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[8]),
        .io_in_control_8_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[8]),
        .io_in_control_8_0_shift(in_input_1_1_payload_Some_0_control_shift[8*5 +: 5]),
        .io_in_control_9_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[9]),
        .io_in_control_9_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[9]),
        .io_in_control_9_0_shift(in_input_1_1_payload_Some_0_control_shift[9*5 +: 5]),
        .io_in_control_10_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[10]),
        .io_in_control_10_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[10]),
        .io_in_control_10_0_shift(in_input_1_1_payload_Some_0_control_shift[10*5 +: 5]),
        .io_in_control_11_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[11]),
        .io_in_control_11_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[11]),
        .io_in_control_11_0_shift(in_input_1_1_payload_Some_0_control_shift[11*5 +: 5]),
        .io_in_control_12_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[12]),
        .io_in_control_12_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[12]),
        .io_in_control_12_0_shift(in_input_1_1_payload_Some_0_control_shift[12*5 +: 5]),
        .io_in_control_13_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[13]),
        .io_in_control_13_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[13]),
        .io_in_control_13_0_shift(in_input_1_1_payload_Some_0_control_shift[13*5 +: 5]),
        .io_in_control_14_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[14]),
        .io_in_control_14_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[14]),
        .io_in_control_14_0_shift(in_input_1_1_payload_Some_0_control_shift[14*5 +: 5]),
        .io_in_control_15_0_dataflow(in_input_1_1_payload_Some_0_control_dataflow_discriminant[15]),
        .io_in_control_15_0_propagate(in_input_1_1_payload_Some_0_control_propagate_discriminant[15]),
        .io_in_control_15_0_shift(in_input_1_1_payload_Some_0_control_shift[15*5 +: 5]),

        .io_in_id_0_0(in_input_1_1_payload_Some_0_id[0*3 +: 3]),
        .io_in_id_1_0(in_input_1_1_payload_Some_0_id[1*3 +: 3]),
        .io_in_id_2_0(in_input_1_1_payload_Some_0_id[2*3 +: 3]),
        .io_in_id_3_0(in_input_1_1_payload_Some_0_id[3*3 +: 3]),
        .io_in_id_4_0(in_input_1_1_payload_Some_0_id[4*3 +: 3]),
        .io_in_id_5_0(in_input_1_1_payload_Some_0_id[5*3 +: 3]),
        .io_in_id_6_0(in_input_1_1_payload_Some_0_id[6*3 +: 3]),
        .io_in_id_7_0(in_input_1_1_payload_Some_0_id[7*3 +: 3]),
        .io_in_id_8_0(in_input_1_1_payload_Some_0_id[8*3 +: 3]),
        .io_in_id_9_0(in_input_1_1_payload_Some_0_id[9*3 +: 3]),
        .io_in_id_10_0(in_input_1_1_payload_Some_0_id[10*3 +: 3]),
        .io_in_id_11_0(in_input_1_1_payload_Some_0_id[11*3 +: 3]),
        .io_in_id_12_0(in_input_1_1_payload_Some_0_id[12*3 +: 3]),
        .io_in_id_13_0(in_input_1_1_payload_Some_0_id[13*3 +: 3]),
        .io_in_id_14_0(in_input_1_1_payload_Some_0_id[14*3 +: 3]),
        .io_in_id_15_0(in_input_1_1_payload_Some_0_id[15*3 +: 3]),

        .io_in_last_0_0(in_input_1_1_payload_Some_0_last[0]),
        .io_in_last_1_0(in_input_1_1_payload_Some_0_last[1]),
        .io_in_last_2_0(in_input_1_1_payload_Some_0_last[2]),
        .io_in_last_3_0(in_input_1_1_payload_Some_0_last[3]),
        .io_in_last_4_0(in_input_1_1_payload_Some_0_last[4]),
        .io_in_last_5_0(in_input_1_1_payload_Some_0_last[5]),
        .io_in_last_6_0(in_input_1_1_payload_Some_0_last[6]),
        .io_in_last_7_0(in_input_1_1_payload_Some_0_last[7]),
        .io_in_last_8_0(in_input_1_1_payload_Some_0_last[8]),
        .io_in_last_9_0(in_input_1_1_payload_Some_0_last[9]),
        .io_in_last_10_0(in_input_1_1_payload_Some_0_last[10]),
        .io_in_last_11_0(in_input_1_1_payload_Some_0_last[11]),
        .io_in_last_12_0(in_input_1_1_payload_Some_0_last[12]),
        .io_in_last_13_0(in_input_1_1_payload_Some_0_last[13]),
        .io_in_last_14_0(in_input_1_1_payload_Some_0_last[14]),
        .io_in_last_15_0(in_input_1_1_payload_Some_0_last[15]),

        .io_in_valid_0_0(in_input_1_1_payload_discriminant[0]),
        .io_in_valid_1_0(in_input_1_1_payload_discriminant[1]),
        .io_in_valid_2_0(in_input_1_1_payload_discriminant[2]),
        .io_in_valid_3_0(in_input_1_1_payload_discriminant[3]),
        .io_in_valid_4_0(in_input_1_1_payload_discriminant[4]),
        .io_in_valid_5_0(in_input_1_1_payload_discriminant[5]),
        .io_in_valid_6_0(in_input_1_1_payload_discriminant[6]),
        .io_in_valid_7_0(in_input_1_1_payload_discriminant[7]),
        .io_in_valid_8_0(in_input_1_1_payload_discriminant[8]),
        .io_in_valid_9_0(in_input_1_1_payload_discriminant[9]),
        .io_in_valid_10_0(in_input_1_1_payload_discriminant[10]),
        .io_in_valid_11_0(in_input_1_1_payload_discriminant[11]),
        .io_in_valid_12_0(in_input_1_1_payload_discriminant[12]),
        .io_in_valid_13_0(in_input_1_1_payload_discriminant[13]),
        .io_in_valid_14_0(in_input_1_1_payload_discriminant[14]),
        .io_in_valid_15_0(in_input_1_1_payload_discriminant[15]),

        .io_out_b_0_0(out_output_1_0_payload_Some_0_b_0[0*20 +: 20]),
        .io_out_b_1_0(out_output_1_0_payload_Some_0_b_0[1*20 +: 20]),
        .io_out_b_2_0(out_output_1_0_payload_Some_0_b_0[2*20 +: 20]),
        .io_out_b_3_0(out_output_1_0_payload_Some_0_b_0[3*20 +: 20]),
        .io_out_b_4_0(out_output_1_0_payload_Some_0_b_0[4*20 +: 20]),
        .io_out_b_5_0(out_output_1_0_payload_Some_0_b_0[5*20 +: 20]),
        .io_out_b_6_0(out_output_1_0_payload_Some_0_b_0[6*20 +: 20]),
        .io_out_b_7_0(out_output_1_0_payload_Some_0_b_0[7*20 +: 20]),
        .io_out_b_8_0(out_output_1_0_payload_Some_0_b_0[8*20 +: 20]),
        .io_out_b_9_0(out_output_1_0_payload_Some_0_b_0[9*20 +: 20]),
        .io_out_b_10_0(out_output_1_0_payload_Some_0_b_0[10*20 +: 20]),
        .io_out_b_11_0(out_output_1_0_payload_Some_0_b_0[11*20 +: 20]),
        .io_out_b_12_0(out_output_1_0_payload_Some_0_b_0[12*20 +: 20]),
        .io_out_b_13_0(out_output_1_0_payload_Some_0_b_0[13*20 +: 20]),
        .io_out_b_14_0(out_output_1_0_payload_Some_0_b_0[14*20 +: 20]),
        .io_out_b_15_0(out_output_1_0_payload_Some_0_b_0[15*20 +: 20]),

        .io_out_c_0_0(out_output_1_0_payload_Some_0_d_0[0*20 +: 20]),
        .io_out_c_1_0(out_output_1_0_payload_Some_0_d_0[1*20 +: 20]),
        .io_out_c_2_0(out_output_1_0_payload_Some_0_d_0[2*20 +: 20]),
        .io_out_c_3_0(out_output_1_0_payload_Some_0_d_0[3*20 +: 20]),
        .io_out_c_4_0(out_output_1_0_payload_Some_0_d_0[4*20 +: 20]),
        .io_out_c_5_0(out_output_1_0_payload_Some_0_d_0[5*20 +: 20]),
        .io_out_c_6_0(out_output_1_0_payload_Some_0_d_0[6*20 +: 20]),
        .io_out_c_7_0(out_output_1_0_payload_Some_0_d_0[7*20 +: 20]),
        .io_out_c_8_0(out_output_1_0_payload_Some_0_d_0[8*20 +: 20]),
        .io_out_c_9_0(out_output_1_0_payload_Some_0_d_0[9*20 +: 20]),
        .io_out_c_10_0(out_output_1_0_payload_Some_0_d_0[10*20 +: 20]),
        .io_out_c_11_0(out_output_1_0_payload_Some_0_d_0[11*20 +: 20]),
        .io_out_c_12_0(out_output_1_0_payload_Some_0_d_0[12*20 +: 20]),
        .io_out_c_13_0(out_output_1_0_payload_Some_0_d_0[13*20 +: 20]),
        .io_out_c_14_0(out_output_1_0_payload_Some_0_d_0[14*20 +: 20]),
        .io_out_c_15_0(out_output_1_0_payload_Some_0_d_0[15*20 +: 20]),

        .io_out_valid_0_0(io_out_valid_0_0),
        .io_out_control_0_0_dataflow(io_out_control_0_0_dataflow),
        .io_out_id_0_0(io_out_id_0_0),
        .io_out_last_0_0(io_out_last_0_0)
    );
    assign out_output_1_0_payload_discriminant[0] = io_out_valid_0_0;
    assign out_output_1_0_payload_discriminant[1] = 1'b1;
    assign out_output_1_0_payload_discriminant[2] = 1'b1;
    assign out_output_1_0_payload_discriminant[3] = 1'b1;
    assign out_output_1_0_payload_discriminant[4] = 1'b1;
    assign out_output_1_0_payload_discriminant[5] = 1'b1;
    assign out_output_1_0_payload_discriminant[6] = 1'b1;
    assign out_output_1_0_payload_discriminant[7] = 1'b1;
    assign out_output_1_0_payload_discriminant[8] = 1'b1;
    assign out_output_1_0_payload_discriminant[9] = 1'b1;
    assign out_output_1_0_payload_discriminant[10] = 1'b1;
    assign out_output_1_0_payload_discriminant[11] = 1'b1;
    assign out_output_1_0_payload_discriminant[12] = 1'b1;
    assign out_output_1_0_payload_discriminant[13] = 1'b1;
    assign out_output_1_0_payload_discriminant[14] = 1'b1;
    assign out_output_1_0_payload_discriminant[15] = 1'b1;

    assign out_output_1_1_payload_discriminant[0] = io_out_valid_0_0;
    assign out_output_1_1_payload_discriminant[1] = 1'b1;
    assign out_output_1_1_payload_discriminant[2] = 1'b1;
    assign out_output_1_1_payload_discriminant[3] = 1'b1;
    assign out_output_1_1_payload_discriminant[4] = 1'b1;
    assign out_output_1_1_payload_discriminant[5] = 1'b1;
    assign out_output_1_1_payload_discriminant[6] = 1'b1;
    assign out_output_1_1_payload_discriminant[7] = 1'b1;
    assign out_output_1_1_payload_discriminant[8] = 1'b1;
    assign out_output_1_1_payload_discriminant[9] = 1'b1;
    assign out_output_1_1_payload_discriminant[10] = 1'b1;
    assign out_output_1_1_payload_discriminant[11] = 1'b1;
    assign out_output_1_1_payload_discriminant[12] = 1'b1;
    assign out_output_1_1_payload_discriminant[13] = 1'b1;
    assign out_output_1_1_payload_discriminant[14] = 1'b1;
    assign out_output_1_1_payload_discriminant[15] = 1'b1;

    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[0] = io_out_control_0_0_dataflow;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[1] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[2] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[3] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[4] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[5] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[6] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[7] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[8] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[9] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[10] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[11] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[12] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[13] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[14] = 1'bx;
    assign out_output_1_1_payload_Some_0_control_dataflow_discriminant[15] = 1'bx;

    assign out_output_1_1_payload_Some_0_id[0*3 +: 3] = io_out_id_0_0;
    assign out_output_1_1_payload_Some_0_id[1*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[2*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[3*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[4*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[5*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[6*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[7*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[8*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[9*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[10*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[11*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[12*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[13*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[14*3 +: 3] = {3{1'bx}};
    assign out_output_1_1_payload_Some_0_id[15*3 +: 3] = {3{1'bx}};

    assign out_output_1_1_payload_Some_0_last[0] = io_out_last_0_0;
    assign out_output_1_1_payload_Some_0_last[1] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[2] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[3] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[4] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[5] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[6] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[7] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[8] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[9] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[10] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[11] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[12] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[13] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[14] = 1'bx;
    assign out_output_1_1_payload_Some_0_last[15] = 1'bx;

endmodule