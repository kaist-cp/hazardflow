// Language: Verilog 2001

`timescale 1ns / 1ps

module fir (
    input  wire             clk,
    input  wire             rst,
    input  wire [8-1:0]     data_in,
    output wire [32-1:0]    data_out
);

// TODO: Implement this module.

initial begin
    $dumpfile("fir.vcd");
    $dumpvars(0, fir);
end

endmodule
