module ReservationStationBlackBoxAdapter (
  input         clock,
                reset,

  input         io_alloc_valid,
  input  [6:0]  io_alloc_bits_cmd_inst_funct,
  input  [4:0]  io_alloc_bits_cmd_inst_rs2,
                io_alloc_bits_cmd_inst_rs1,
  input         io_alloc_bits_cmd_inst_xd,
                io_alloc_bits_cmd_inst_xs1,
                io_alloc_bits_cmd_inst_xs2,
  input  [4:0]  io_alloc_bits_cmd_inst_rd,
  input  [6:0]  io_alloc_bits_cmd_inst_opcode,
  input  [63:0] io_alloc_bits_cmd_rs1,
                io_alloc_bits_cmd_rs2,
  input         io_alloc_bits_cmd_status_debug,
                io_alloc_bits_cmd_status_cease,
                io_alloc_bits_cmd_status_wfi,
  input  [31:0] io_alloc_bits_cmd_status_isa,
  input  [1:0]  io_alloc_bits_cmd_status_dprv,
  input         io_alloc_bits_cmd_status_dv,
  input  [1:0]  io_alloc_bits_cmd_status_prv,
  input         io_alloc_bits_cmd_status_v,
                io_alloc_bits_cmd_status_sd,
  input  [22:0] io_alloc_bits_cmd_status_zero2,
  input         io_alloc_bits_cmd_status_mpv,
                io_alloc_bits_cmd_status_gva,
                io_alloc_bits_cmd_status_mbe,
                io_alloc_bits_cmd_status_sbe,
  input  [1:0]  io_alloc_bits_cmd_status_sxl,
                io_alloc_bits_cmd_status_uxl,
  input         io_alloc_bits_cmd_status_sd_rv32,
  input  [7:0]  io_alloc_bits_cmd_status_zero1,
  input         io_alloc_bits_cmd_status_tsr,
                io_alloc_bits_cmd_status_tw,
                io_alloc_bits_cmd_status_tvm,
                io_alloc_bits_cmd_status_mxr,
                io_alloc_bits_cmd_status_sum,
                io_alloc_bits_cmd_status_mprv,
  input  [1:0]  io_alloc_bits_cmd_status_xs,
                io_alloc_bits_cmd_status_fs,
                io_alloc_bits_cmd_status_mpp,
                io_alloc_bits_cmd_status_vs,
  input         io_alloc_bits_cmd_status_spp,
                io_alloc_bits_cmd_status_mpie,
                io_alloc_bits_cmd_status_ube,
                io_alloc_bits_cmd_status_spie,
                io_alloc_bits_cmd_status_upie,
                io_alloc_bits_cmd_status_mie,
                io_alloc_bits_cmd_status_hie,
                io_alloc_bits_cmd_status_sie,
                io_alloc_bits_cmd_status_uie,
                io_alloc_bits_from_matmul_fsm,
                io_alloc_bits_from_conv_fsm,
  output        io_alloc_ready,

  input         io_completed_valid,
  input  [5:0]  io_completed_bits,

  input         io_issue_ld_ready,
  output        io_issue_ld_valid,
  output [6:0]  io_issue_ld_cmd_cmd_inst_funct,
  output [4:0]  io_issue_ld_cmd_cmd_inst_rs2,
                io_issue_ld_cmd_cmd_inst_rs1,
  output        io_issue_ld_cmd_cmd_inst_xd,
                io_issue_ld_cmd_cmd_inst_xs1,
                io_issue_ld_cmd_cmd_inst_xs2,
  output [4:0]  io_issue_ld_cmd_cmd_inst_rd,
  output [6:0]  io_issue_ld_cmd_cmd_inst_opcode,
  output [63:0] io_issue_ld_cmd_cmd_rs1,
                io_issue_ld_cmd_cmd_rs2,
  output        io_issue_ld_cmd_cmd_status_debug,
                io_issue_ld_cmd_cmd_status_cease,
                io_issue_ld_cmd_cmd_status_wfi,
  output [31:0] io_issue_ld_cmd_cmd_status_isa,
  output [1:0]  io_issue_ld_cmd_cmd_status_dprv,
  output        io_issue_ld_cmd_cmd_status_dv,
  output [1:0]  io_issue_ld_cmd_cmd_status_prv,
  output        io_issue_ld_cmd_cmd_status_v,
                io_issue_ld_cmd_cmd_status_sd,
  output [22:0] io_issue_ld_cmd_cmd_status_zero2,
  output        io_issue_ld_cmd_cmd_status_mpv,
                io_issue_ld_cmd_cmd_status_gva,
                io_issue_ld_cmd_cmd_status_mbe,
                io_issue_ld_cmd_cmd_status_sbe,
  output [1:0]  io_issue_ld_cmd_cmd_status_sxl,
                io_issue_ld_cmd_cmd_status_uxl,
  output        io_issue_ld_cmd_cmd_status_sd_rv32,
  output [7:0]  io_issue_ld_cmd_cmd_status_zero1,
  output        io_issue_ld_cmd_cmd_status_tsr,
                io_issue_ld_cmd_cmd_status_tw,
                io_issue_ld_cmd_cmd_status_tvm,
                io_issue_ld_cmd_cmd_status_mxr,
                io_issue_ld_cmd_cmd_status_sum,
                io_issue_ld_cmd_cmd_status_mprv,
  output [1:0]  io_issue_ld_cmd_cmd_status_xs,
                io_issue_ld_cmd_cmd_status_fs,
                io_issue_ld_cmd_cmd_status_mpp,
                io_issue_ld_cmd_cmd_status_vs,
  output        io_issue_ld_cmd_cmd_status_spp,
                io_issue_ld_cmd_cmd_status_mpie,
                io_issue_ld_cmd_cmd_status_ube,
                io_issue_ld_cmd_cmd_status_spie,
                io_issue_ld_cmd_cmd_status_upie,
                io_issue_ld_cmd_cmd_status_mie,
                io_issue_ld_cmd_cmd_status_hie,
                io_issue_ld_cmd_cmd_status_sie,
                io_issue_ld_cmd_cmd_status_uie,
                io_issue_ld_cmd_from_matmul_fsm,
                io_issue_ld_cmd_from_conv_fsm,
  output [5:0]  io_issue_ld_rob_id,

  input         io_issue_st_ready,
  output        io_issue_st_valid,
  output [6:0]  io_issue_st_cmd_cmd_inst_funct,
  output [4:0]  io_issue_st_cmd_cmd_inst_rs2,
                io_issue_st_cmd_cmd_inst_rs1,
  output        io_issue_st_cmd_cmd_inst_xd,
                io_issue_st_cmd_cmd_inst_xs1,
                io_issue_st_cmd_cmd_inst_xs2,
  output [4:0]  io_issue_st_cmd_cmd_inst_rd,
  output [6:0]  io_issue_st_cmd_cmd_inst_opcode,
  output [63:0] io_issue_st_cmd_cmd_rs1,
                io_issue_st_cmd_cmd_rs2,
  output        io_issue_st_cmd_cmd_status_debug,
                io_issue_st_cmd_cmd_status_cease,
                io_issue_st_cmd_cmd_status_wfi,
  output [31:0] io_issue_st_cmd_cmd_status_isa,
  output [1:0]  io_issue_st_cmd_cmd_status_dprv,
  output        io_issue_st_cmd_cmd_status_dv,
  output [1:0]  io_issue_st_cmd_cmd_status_prv,
  output        io_issue_st_cmd_cmd_status_v,
                io_issue_st_cmd_cmd_status_sd,
  output [22:0] io_issue_st_cmd_cmd_status_zero2,
  output        io_issue_st_cmd_cmd_status_mpv,
                io_issue_st_cmd_cmd_status_gva,
                io_issue_st_cmd_cmd_status_mbe,
                io_issue_st_cmd_cmd_status_sbe,
  output [1:0]  io_issue_st_cmd_cmd_status_sxl,
                io_issue_st_cmd_cmd_status_uxl,
  output        io_issue_st_cmd_cmd_status_sd_rv32,
  output [7:0]  io_issue_st_cmd_cmd_status_zero1,
  output        io_issue_st_cmd_cmd_status_tsr,
                io_issue_st_cmd_cmd_status_tw,
                io_issue_st_cmd_cmd_status_tvm,
                io_issue_st_cmd_cmd_status_mxr,
                io_issue_st_cmd_cmd_status_sum,
                io_issue_st_cmd_cmd_status_mprv,
  output [1:0]  io_issue_st_cmd_cmd_status_xs,
                io_issue_st_cmd_cmd_status_fs,
                io_issue_st_cmd_cmd_status_mpp,
                io_issue_st_cmd_cmd_status_vs,
  output        io_issue_st_cmd_cmd_status_spp,
                io_issue_st_cmd_cmd_status_mpie,
                io_issue_st_cmd_cmd_status_ube,
                io_issue_st_cmd_cmd_status_spie,
                io_issue_st_cmd_cmd_status_upie,
                io_issue_st_cmd_cmd_status_mie,
                io_issue_st_cmd_cmd_status_hie,
                io_issue_st_cmd_cmd_status_sie,
                io_issue_st_cmd_cmd_status_uie,
                io_issue_st_cmd_from_matmul_fsm,
                io_issue_st_cmd_from_conv_fsm,
  output [5:0]  io_issue_st_rob_id,

  input         io_issue_ex_ready,
  output        io_issue_ex_valid,
  output [6:0]  io_issue_ex_cmd_cmd_inst_funct,
  output [63:0] io_issue_ex_cmd_cmd_rs1,
                io_issue_ex_cmd_cmd_rs2,
  output [5:0]  io_issue_ex_rob_id,

  output [1:0]  io_conv_ld_completed,
                io_conv_ex_completed,
                io_conv_st_completed,

  output [1:0]  io_matmul_ld_completed,
                io_matmul_ex_completed,
                io_matmul_st_completed,

  output        io_busy
);

reservation_station_top reservation_station(
  .clk(clock),
  .rst(reset),

  .in_input_0_payload_discriminant(io_alloc_valid),
  .in_input_0_payload_Some_0_cmd_inst_funct_discriminant(io_alloc_bits_cmd_inst_funct),
  .in_input_0_payload_Some_0_cmd_inst_rs2(io_alloc_bits_cmd_inst_rs2),
  .in_input_0_payload_Some_0_cmd_inst_rs1(io_alloc_bits_cmd_inst_rs1),
  .in_input_0_payload_Some_0_cmd_inst_xd(io_alloc_bits_cmd_inst_xd),
  .in_input_0_payload_Some_0_cmd_inst_xs1(io_alloc_bits_cmd_inst_xs1),
  .in_input_0_payload_Some_0_cmd_inst_xs2(io_alloc_bits_cmd_inst_xs2),
  .in_input_0_payload_Some_0_cmd_inst_rd(io_alloc_bits_cmd_inst_rd),
  .in_input_0_payload_Some_0_cmd_inst_opcode(io_alloc_bits_cmd_inst_opcode),
  .in_input_0_payload_Some_0_cmd_rs1(io_alloc_bits_cmd_rs1),
  .in_input_0_payload_Some_0_cmd_rs2(io_alloc_bits_cmd_rs2),
  .in_input_0_payload_Some_0_cmd_status_debug(io_alloc_bits_cmd_status_debug),
  .in_input_0_payload_Some_0_cmd_status_cease(io_alloc_bits_cmd_status_cease),
  .in_input_0_payload_Some_0_cmd_status_wfi(io_alloc_bits_cmd_status_wfi),
  .in_input_0_payload_Some_0_cmd_status_isa(io_alloc_bits_cmd_status_isa),
  .in_input_0_payload_Some_0_cmd_status_dprv(io_alloc_bits_cmd_status_dprv),
  .in_input_0_payload_Some_0_cmd_status_dv(io_alloc_bits_cmd_status_dv),
  .in_input_0_payload_Some_0_cmd_status_prv(io_alloc_bits_cmd_status_prv),
  .in_input_0_payload_Some_0_cmd_status_v(io_alloc_bits_cmd_status_v),
  .in_input_0_payload_Some_0_cmd_status_sd(io_alloc_bits_cmd_status_sd),
  .in_input_0_payload_Some_0_cmd_status_zero2(io_alloc_bits_cmd_status_zero2),
  .in_input_0_payload_Some_0_cmd_status_mpv(io_alloc_bits_cmd_status_mpv),
  .in_input_0_payload_Some_0_cmd_status_gva(io_alloc_bits_cmd_status_gva),
  .in_input_0_payload_Some_0_cmd_status_mbe(io_alloc_bits_cmd_status_mbe),
  .in_input_0_payload_Some_0_cmd_status_sbe(io_alloc_bits_cmd_status_sbe),
  .in_input_0_payload_Some_0_cmd_status_sxl(io_alloc_bits_cmd_status_sxl),
  .in_input_0_payload_Some_0_cmd_status_uxl(io_alloc_bits_cmd_status_uxl),
  .in_input_0_payload_Some_0_cmd_status_sd_rv32(io_alloc_bits_cmd_status_sd_rv32),
  .in_input_0_payload_Some_0_cmd_status_zero1(io_alloc_bits_cmd_status_zero1),
  .in_input_0_payload_Some_0_cmd_status_tsr(io_alloc_bits_cmd_status_tsr),
  .in_input_0_payload_Some_0_cmd_status_tw(io_alloc_bits_cmd_status_tw),
  .in_input_0_payload_Some_0_cmd_status_tvm(io_alloc_bits_cmd_status_tvm),
  .in_input_0_payload_Some_0_cmd_status_mxr(io_alloc_bits_cmd_status_mxr),
  .in_input_0_payload_Some_0_cmd_status_sum(io_alloc_bits_cmd_status_sum),
  .in_input_0_payload_Some_0_cmd_status_mprv(io_alloc_bits_cmd_status_mprv),
  .in_input_0_payload_Some_0_cmd_status_xs(io_alloc_bits_cmd_status_xs),
  .in_input_0_payload_Some_0_cmd_status_fs(io_alloc_bits_cmd_status_fs),
  .in_input_0_payload_Some_0_cmd_status_mpp(io_alloc_bits_cmd_status_mpp),
  .in_input_0_payload_Some_0_cmd_status_vs(io_alloc_bits_cmd_status_vs),
  .in_input_0_payload_Some_0_cmd_status_spp(io_alloc_bits_cmd_status_spp),
  .in_input_0_payload_Some_0_cmd_status_mpie(io_alloc_bits_cmd_status_mpie),
  .in_input_0_payload_Some_0_cmd_status_ube(io_alloc_bits_cmd_status_ube),
  .in_input_0_payload_Some_0_cmd_status_spie(io_alloc_bits_cmd_status_spie),
  .in_input_0_payload_Some_0_cmd_status_upie(io_alloc_bits_cmd_status_upie),
  .in_input_0_payload_Some_0_cmd_status_mie(io_alloc_bits_cmd_status_mie),
  .in_input_0_payload_Some_0_cmd_status_hie(io_alloc_bits_cmd_status_hie),
  .in_input_0_payload_Some_0_cmd_status_sie(io_alloc_bits_cmd_status_sie),
  .in_input_0_payload_Some_0_cmd_status_uie(io_alloc_bits_cmd_status_uie),
  .in_input_0_payload_Some_0_rob_id_discriminant(),
  .in_input_0_payload_Some_0_rob_id_Some_0(),
  .in_input_0_payload_Some_0_from_matmul_fsm(io_alloc_bits_from_matmul_fsm),
  .in_input_0_payload_Some_0_from_conv_fsm(io_alloc_bits_from_conv_fsm),
  .in_input_0_resolver_ready(io_alloc_ready),

  .in_input_1_payload_discriminant(io_completed_valid),
  .in_input_1_payload_Some_0(io_completed_bits),

  .out_output_0_ld_resolver_ready(io_issue_ld_ready),
  .out_output_0_ld_payload_discriminant(io_issue_ld_valid),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_funct_discriminant(io_issue_ld_cmd_cmd_inst_funct),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_rs2(io_issue_ld_cmd_cmd_inst_rs2),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_rs1(io_issue_ld_cmd_cmd_inst_rs1),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_xd(io_issue_ld_cmd_cmd_inst_xd),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_xs1(io_issue_ld_cmd_cmd_inst_xs1),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_xs2(io_issue_ld_cmd_cmd_inst_xs2),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_rd(io_issue_ld_cmd_cmd_inst_rd),
  .out_output_0_ld_payload_Some_0_cmd_cmd_inst_opcode(io_issue_ld_cmd_cmd_inst_opcode),
  .out_output_0_ld_payload_Some_0_cmd_cmd_rs1(io_issue_ld_cmd_cmd_rs1),
  .out_output_0_ld_payload_Some_0_cmd_cmd_rs2(io_issue_ld_cmd_cmd_rs2),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_debug(io_issue_ld_cmd_cmd_status_debug),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_cease(io_issue_ld_cmd_cmd_status_cease),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_wfi(io_issue_ld_cmd_cmd_status_wfi),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_isa(io_issue_ld_cmd_cmd_status_isa),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_dprv(io_issue_ld_cmd_cmd_status_dprv),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_dv(io_issue_ld_cmd_cmd_status_dv),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_prv(io_issue_ld_cmd_cmd_status_prv),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_v(io_issue_ld_cmd_cmd_status_v),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sd(io_issue_ld_cmd_cmd_status_sd),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_zero2(io_issue_ld_cmd_cmd_status_zero2),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mpv(io_issue_ld_cmd_cmd_status_mpv),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_gva(io_issue_ld_cmd_cmd_status_gva),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mbe(io_issue_ld_cmd_cmd_status_mbe),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sbe(io_issue_ld_cmd_cmd_status_sbe),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sxl(io_issue_ld_cmd_cmd_status_sxl),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_uxl(io_issue_ld_cmd_cmd_status_uxl),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sd_rv32(io_issue_ld_cmd_cmd_status_sd_rv32),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_zero1(io_issue_ld_cmd_cmd_status_zero1),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_tsr(io_issue_ld_cmd_cmd_status_tsr),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_tw(io_issue_ld_cmd_cmd_status_tw),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_tvm(io_issue_ld_cmd_cmd_status_tvm),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mxr(io_issue_ld_cmd_cmd_status_mxr),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sum(io_issue_ld_cmd_cmd_status_sum),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mprv(io_issue_ld_cmd_cmd_status_mprv),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_xs(io_issue_ld_cmd_cmd_status_xs),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_fs(io_issue_ld_cmd_cmd_status_fs),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mpp(io_issue_ld_cmd_cmd_status_mpp),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_vs(io_issue_ld_cmd_cmd_status_vs),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_spp(io_issue_ld_cmd_cmd_status_spp),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mpie(io_issue_ld_cmd_cmd_status_mpie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_ube(io_issue_ld_cmd_cmd_status_ube),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_spie(io_issue_ld_cmd_cmd_status_spie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_upie(io_issue_ld_cmd_cmd_status_upie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_mie(io_issue_ld_cmd_cmd_status_mie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_hie(io_issue_ld_cmd_cmd_status_hie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_sie(io_issue_ld_cmd_cmd_status_sie),
  .out_output_0_ld_payload_Some_0_cmd_cmd_status_uie(io_issue_ld_cmd_cmd_status_uie),
  .out_output_0_ld_payload_Some_0_cmd_rob_id_discriminant(),
  .out_output_0_ld_payload_Some_0_cmd_rob_id_Some_0(),
  .out_output_0_ld_payload_Some_0_cmd_from_matmul_fsm(io_issue_ld_cmd_from_matmul_fsm),
  .out_output_0_ld_payload_Some_0_cmd_from_conv_fsm(io_issue_ld_cmd_from_conv_fsm),
  .out_output_0_ld_payload_Some_0_rob_id(io_issue_ld_rob_id),

  .out_output_0_st_resolver_ready(io_issue_st_ready),
  .out_output_0_st_payload_discriminant(io_issue_st_valid),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_funct_discriminant(io_issue_st_cmd_cmd_inst_funct),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_rs2(io_issue_st_cmd_cmd_inst_rs2),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_rs1(io_issue_st_cmd_cmd_inst_rs1),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_xd(io_issue_st_cmd_cmd_inst_xd),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_xs1(io_issue_st_cmd_cmd_inst_xs1),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_xs2(io_issue_st_cmd_cmd_inst_xs2),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_rd(io_issue_st_cmd_cmd_inst_rd),
  .out_output_0_st_payload_Some_0_cmd_cmd_inst_opcode(io_issue_st_cmd_cmd_inst_opcode),
  .out_output_0_st_payload_Some_0_cmd_cmd_rs1(io_issue_st_cmd_cmd_rs1),
  .out_output_0_st_payload_Some_0_cmd_cmd_rs2(io_issue_st_cmd_cmd_rs2),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_debug(io_issue_st_cmd_cmd_status_debug),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_cease(io_issue_st_cmd_cmd_status_cease),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_wfi(io_issue_st_cmd_cmd_status_wfi),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_isa(io_issue_st_cmd_cmd_status_isa),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_dprv(io_issue_st_cmd_cmd_status_dprv),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_dv(io_issue_st_cmd_cmd_status_dv),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_prv(io_issue_st_cmd_cmd_status_prv),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_v(io_issue_st_cmd_cmd_status_v),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sd(io_issue_st_cmd_cmd_status_sd),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_zero2(io_issue_st_cmd_cmd_status_zero2),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mpv(io_issue_st_cmd_cmd_status_mpv),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_gva(io_issue_st_cmd_cmd_status_gva),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mbe(io_issue_st_cmd_cmd_status_mbe),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sbe(io_issue_st_cmd_cmd_status_sbe),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sxl(io_issue_st_cmd_cmd_status_sxl),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_uxl(io_issue_st_cmd_cmd_status_uxl),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sd_rv32(io_issue_st_cmd_cmd_status_sd_rv32),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_zero1(io_issue_st_cmd_cmd_status_zero1),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_tsr(io_issue_st_cmd_cmd_status_tsr),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_tw(io_issue_st_cmd_cmd_status_tw),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_tvm(io_issue_st_cmd_cmd_status_tvm),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mxr(io_issue_st_cmd_cmd_status_mxr),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sum(io_issue_st_cmd_cmd_status_sum),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mprv(io_issue_st_cmd_cmd_status_mprv),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_xs(io_issue_st_cmd_cmd_status_xs),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_fs(io_issue_st_cmd_cmd_status_fs),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mpp(io_issue_st_cmd_cmd_status_mpp),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_vs(io_issue_st_cmd_cmd_status_vs),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_spp(io_issue_st_cmd_cmd_status_spp),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mpie(io_issue_st_cmd_cmd_status_mpie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_ube(io_issue_st_cmd_cmd_status_ube),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_spie(io_issue_st_cmd_cmd_status_spie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_upie(io_issue_st_cmd_cmd_status_upie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_mie(io_issue_st_cmd_cmd_status_mie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_hie(io_issue_st_cmd_cmd_status_hie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_sie(io_issue_st_cmd_cmd_status_sie),
  .out_output_0_st_payload_Some_0_cmd_cmd_status_uie(io_issue_st_cmd_cmd_status_uie),
  .out_output_0_st_payload_Some_0_cmd_rob_id_discriminant(),
  .out_output_0_st_payload_Some_0_cmd_rob_id_Some_0(),
  .out_output_0_st_payload_Some_0_cmd_from_matmul_fsm(io_issue_st_cmd_from_matmul_fsm),
  .out_output_0_st_payload_Some_0_cmd_from_conv_fsm(io_issue_st_cmd_from_conv_fsm),
  .out_output_0_st_payload_Some_0_rob_id(io_issue_st_rob_id),

  .out_output_0_ex_resolver_ready(io_issue_ex_ready),
  .out_output_0_ex_payload_discriminant(io_issue_ex_valid),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_funct_discriminant(io_issue_ex_cmd_cmd_inst_funct),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_rs2(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_rs1(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_xd(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_xs1(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_xs2(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_rd(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_inst_opcode(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_rs1(io_issue_ex_cmd_cmd_rs1),
  .out_output_0_ex_payload_Some_0_cmd_cmd_rs2(io_issue_ex_cmd_cmd_rs2),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_debug(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_cease(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_wfi(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_isa(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_dprv(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_dv(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_prv(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_v(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sd(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_zero2(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mpv(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_gva(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mbe(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sbe(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sxl(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_uxl(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sd_rv32(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_zero1(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_tsr(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_tw(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_tvm(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mxr(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sum(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mprv(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_xs(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_fs(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mpp(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_vs(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_spp(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mpie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_ube(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_spie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_upie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_mie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_hie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_sie(),
  .out_output_0_ex_payload_Some_0_cmd_cmd_status_uie(),
  .out_output_0_ex_payload_Some_0_cmd_rob_id_discriminant(),
  .out_output_0_ex_payload_Some_0_cmd_rob_id_Some_0(),
  .out_output_0_ex_payload_Some_0_cmd_from_matmul_fsm(),
  .out_output_0_ex_payload_Some_0_cmd_from_conv_fsm(),
  .out_output_0_ex_payload_Some_0_rob_id(io_issue_ex_rob_id),

  .out_output_1_conv_ld_payload_discriminant(),
  .out_output_1_conv_ld_payload_Some_0(io_conv_ld_completed),
  .out_output_1_conv_ex_payload_discriminant(),
  .out_output_1_conv_ex_payload_Some_0(io_conv_ex_completed),
  .out_output_1_conv_st_payload_discriminant(),
  .out_output_1_conv_st_payload_Some_0(io_conv_st_completed),
  .out_output_1_matmul_ld_payload_discriminant(),
  .out_output_1_matmul_ld_payload_Some_0(io_matmul_ld_completed),
  .out_output_1_matmul_ex_payload_discriminant(),
  .out_output_1_matmul_ex_payload_Some_0(io_matmul_ex_completed),
  .out_output_1_matmul_st_payload_discriminant(),
  .out_output_1_matmul_st_payload_Some_0(io_matmul_st_completed),

  .out_output_2_payload_discriminant(),
  .out_output_2_payload_Some_0(io_busy)
);

endmodule
