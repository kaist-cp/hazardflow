module MeshWithDelaysWrapper(
    input wire clk,
    input wire rst,
    input wire in_input_0_0_payload_discriminant,
    input wire [128-1:0] in_input_0_0_payload_Some_0,
    output wire in_input_0_0_resolver_ready,
    input wire in_input_0_1_payload_discriminant,
    input wire [128-1:0] in_input_0_1_payload_Some_0,
    output wire in_input_0_1_resolver_ready,
    input wire in_input_0_2_payload_discriminant,
    input wire [128-1:0] in_input_0_2_payload_Some_0,
    output wire in_input_0_2_resolver_ready,
    input wire in_input_0_3_payload_discriminant,
    input wire in_input_0_3_payload_Some_0_pe_control_dataflow_discriminant,
    input wire in_input_0_3_payload_Some_0_pe_control_propagate_discriminant,
    input wire [5-1:0] in_input_0_3_payload_Some_0_pe_control_shift,
    input wire in_input_0_3_payload_Some_0_transpose_a,
    input wire in_input_0_3_payload_Some_0_transpose_bd,
    input wire [5-1:0] in_input_0_3_payload_Some_0_total_rows,
    input wire in_input_0_3_payload_Some_0_tag_rob_id_discriminant,
    input wire [6-1:0] in_input_0_3_payload_Some_0_tag_rob_id_Some_0,
    input wire in_input_0_3_payload_Some_0_tag_addr_is_acc_addr,
    input wire in_input_0_3_payload_Some_0_tag_addr_accumulate,
    input wire in_input_0_3_payload_Some_0_tag_addr_read_full_acc_row,
    input wire [3-1:0] in_input_0_3_payload_Some_0_tag_addr_norm_cmd,
    input wire [11-1:0] in_input_0_3_payload_Some_0_tag_addr_garbage,
    input wire in_input_0_3_payload_Some_0_tag_addr_is_garbage,
    input wire [14-1:0] in_input_0_3_payload_Some_0_tag_addr_data,
    input wire [5-1:0] in_input_0_3_payload_Some_0_tag_rows,
    input wire [5-1:0] in_input_0_3_payload_Some_0_tag_cols,
    input wire [2-1:0] in_input_0_3_payload_Some_0_flush,

    output wire in_input_0_3_resolver_ready,
    output wire [6-1:0] in_input_0_3_resolver_inner_rob_id_discriminant,
    output wire [36-1:0] in_input_0_3_resolver_inner_rob_id_Some_0,
    output wire [6-1:0] in_input_0_3_resolver_inner_addr_is_acc_addr,
    output wire [6-1:0] in_input_0_3_resolver_inner_addr_accumulate,
    output wire [6-1:0] in_input_0_3_resolver_inner_addr_read_full_acc_row,
    output wire [18-1:0] in_input_0_3_resolver_inner_addr_norm_cmd,
    output wire [66-1:0] in_input_0_3_resolver_inner_addr_garbage,
    output wire [6-1:0] in_input_0_3_resolver_inner_addr_is_garbage,
    output wire [84-1:0] in_input_0_3_resolver_inner_addr_data,
    output wire [30-1:0] in_input_0_3_resolver_inner_rows,
    output wire [30-1:0] in_input_0_3_resolver_inner_cols,
    
    output wire out_output_payload_discriminant,
    output wire [5-1:0] out_output_payload_Some_0_total_rows,
    output wire out_output_payload_Some_0_tag_rob_id_discriminant,
    output wire [6-1:0] out_output_payload_Some_0_tag_rob_id_Some_0,
    output wire out_output_payload_Some_0_tag_addr_is_acc_addr,
    output wire out_output_payload_Some_0_tag_addr_accumulate,
    output wire out_output_payload_Some_0_tag_addr_read_full_acc_row,
    output wire [3-1:0] out_output_payload_Some_0_tag_addr_norm_cmd,
    output wire [11-1:0] out_output_payload_Some_0_tag_addr_garbage,
    output wire out_output_payload_Some_0_tag_addr_is_garbage,
    output wire [14-1:0] out_output_payload_Some_0_tag_addr_data,
    output wire [5-1:0] out_output_payload_Some_0_tag_rows,
    output wire [5-1:0] out_output_payload_Some_0_tag_cols,
    output wire out_output_payload_Some_0_last,
    output wire [320-1:0] out_output_payload_Some_0_data
);

MeshWithDelays mesh_with_delays(
    .clock(clk),
    .reset(rst),
    .io_a_valid(in_input_0_0_payload_discriminant),
    .io_a_bits_0_0(in_input_0_0_payload_Some_0[0*8 +: 8]),
    .io_a_bits_1_0(in_input_0_0_payload_Some_0[1*8 +: 8]),
    .io_a_bits_2_0(in_input_0_0_payload_Some_0[2*8 +: 8]),
    .io_a_bits_3_0(in_input_0_0_payload_Some_0[3*8 +: 8]),
    .io_a_bits_4_0(in_input_0_0_payload_Some_0[4*8 +: 8]),
    .io_a_bits_5_0(in_input_0_0_payload_Some_0[5*8 +: 8]),
    .io_a_bits_6_0(in_input_0_0_payload_Some_0[6*8 +: 8]),
    .io_a_bits_7_0(in_input_0_0_payload_Some_0[7*8 +: 8]),
    .io_a_bits_8_0(in_input_0_0_payload_Some_0[8*8 +: 8]),
    .io_a_bits_9_0(in_input_0_0_payload_Some_0[9*8 +: 8]),
    .io_a_bits_10_0(in_input_0_0_payload_Some_0[10*8 +: 8]),
    .io_a_bits_11_0(in_input_0_0_payload_Some_0[11*8 +: 8]),
    .io_a_bits_12_0(in_input_0_0_payload_Some_0[12*8 +: 8]),
    .io_a_bits_13_0(in_input_0_0_payload_Some_0[13*8 +: 8]),
    .io_a_bits_14_0(in_input_0_0_payload_Some_0[14*8 +: 8]),
    .io_a_bits_15_0(in_input_0_0_payload_Some_0[15*8 +: 8]),
    .io_b_valid(in_input_0_1_payload_discriminant),
    .io_b_bits_0_0(in_input_0_1_payload_Some_0[0*8 +: 8]),
    .io_b_bits_1_0(in_input_0_1_payload_Some_0[1*8 +: 8]),
    .io_b_bits_2_0(in_input_0_1_payload_Some_0[2*8 +: 8]),
    .io_b_bits_3_0(in_input_0_1_payload_Some_0[3*8 +: 8]),
    .io_b_bits_4_0(in_input_0_1_payload_Some_0[4*8 +: 8]),
    .io_b_bits_5_0(in_input_0_1_payload_Some_0[5*8 +: 8]),
    .io_b_bits_6_0(in_input_0_1_payload_Some_0[6*8 +: 8]),
    .io_b_bits_7_0(in_input_0_1_payload_Some_0[7*8 +: 8]),
    .io_b_bits_8_0(in_input_0_1_payload_Some_0[8*8 +: 8]),
    .io_b_bits_9_0(in_input_0_1_payload_Some_0[9*8 +: 8]),
    .io_b_bits_10_0(in_input_0_1_payload_Some_0[10*8 +: 8]),
    .io_b_bits_11_0(in_input_0_1_payload_Some_0[11*8 +: 8]),
    .io_b_bits_12_0(in_input_0_1_payload_Some_0[12*8 +: 8]),
    .io_b_bits_13_0(in_input_0_1_payload_Some_0[13*8 +: 8]),
    .io_b_bits_14_0(in_input_0_1_payload_Some_0[14*8 +: 8]),
    .io_b_bits_15_0(in_input_0_1_payload_Some_0[15*8 +: 8]),
    .io_d_valid(in_input_0_2_payload_discriminant),
    .io_d_bits_0_0(in_input_0_2_payload_Some_0[0*8 +: 8]),
    .io_d_bits_1_0(in_input_0_2_payload_Some_0[1*8 +: 8]),
    .io_d_bits_2_0(in_input_0_2_payload_Some_0[2*8 +: 8]),
    .io_d_bits_3_0(in_input_0_2_payload_Some_0[3*8 +: 8]),
    .io_d_bits_4_0(in_input_0_2_payload_Some_0[4*8 +: 8]),
    .io_d_bits_5_0(in_input_0_2_payload_Some_0[5*8 +: 8]),
    .io_d_bits_6_0(in_input_0_2_payload_Some_0[6*8 +: 8]),
    .io_d_bits_7_0(in_input_0_2_payload_Some_0[7*8 +: 8]),
    .io_d_bits_8_0(in_input_0_2_payload_Some_0[8*8 +: 8]),
    .io_d_bits_9_0(in_input_0_2_payload_Some_0[9*8 +: 8]),
    .io_d_bits_10_0(in_input_0_2_payload_Some_0[10*8 +: 8]),
    .io_d_bits_11_0(in_input_0_2_payload_Some_0[11*8 +: 8]),
    .io_d_bits_12_0(in_input_0_2_payload_Some_0[12*8 +: 8]),
    .io_d_bits_13_0(in_input_0_2_payload_Some_0[13*8 +: 8]),
    .io_d_bits_14_0(in_input_0_2_payload_Some_0[14*8 +: 8]),
    .io_d_bits_15_0(in_input_0_2_payload_Some_0[15*8 +: 8]),
    .io_req_valid(in_input_0_3_payload_discriminant),
    .io_req_bits_tag_rob_id_valid(in_input_0_3_payload_Some_0_tag_rob_id_discriminant),
    .io_req_bits_tag_rob_id_bits(in_input_0_3_payload_Some_0_tag_rob_id_Some_0),
    .io_req_bits_tag_addr_is_acc_addr(in_input_0_3_payload_Some_0_tag_addr_is_acc_addr),
    .io_req_bits_tag_addr_accumulate(in_input_0_3_payload_Some_0_tag_addr_accumulate),
    .io_req_bits_tag_addr_read_full_acc_row(in_input_0_3_payload_Some_0_tag_addr_read_full_acc_row),
    .io_req_bits_tag_addr_garbage_bit(in_input_0_3_payload_Some_0_tag_addr_is_garbage),
    .io_req_bits_tag_addr_data(in_input_0_3_payload_Some_0_tag_addr_data),
    .io_req_bits_tag_rows(in_input_0_3_payload_Some_0_tag_rows),
    .io_req_bits_tag_cols(in_input_0_3_payload_Some_0_tag_cols),
    .io_req_bits_pe_control_dataflow(in_input_0_3_payload_Some_0_pe_control_dataflow_discriminant),
    .io_req_bits_pe_control_propagate(in_input_0_3_payload_Some_0_pe_control_propagate_discriminant),
    .io_req_bits_pe_control_shift(in_input_0_3_payload_Some_0_pe_control_shift),
    .io_req_bits_a_transpose(in_input_0_3_payload_Some_0_transpose_a),
    .io_req_bits_bd_transpose(in_input_0_3_payload_Some_0_transpose_bd),
    .io_req_bits_total_rows(in_input_0_3_payload_Some_0_total_rows),
    .io_req_bits_flush(in_input_0_3_payload_Some_0_flush),
    .io_a_ready(in_input_0_0_resolver_ready),
    .io_b_ready(in_input_0_1_resolver_ready),
    .io_d_ready(in_input_0_2_resolver_ready),
    .io_req_ready(in_input_0_3_resolver_ready),
    .io_resp_valid(out_output_payload_discriminant),
    .io_resp_bits_tag_rob_id_valid(out_output_payload_Some_0_tag_rob_id_discriminant),
    .io_resp_bits_tag_rob_id_bits(out_output_payload_Some_0_tag_rob_id_Some_0),
    .io_resp_bits_tag_addr_is_acc_addr(out_output_payload_Some_0_tag_addr_is_acc_addr),
    .io_resp_bits_tag_addr_accumulate(out_output_payload_Some_0_tag_addr_accumulate),
    .io_resp_bits_tag_addr_read_full_acc_row(out_output_payload_Some_0_tag_addr_read_full_acc_row),
    .io_resp_bits_tag_addr_garbage_bit(out_output_payload_Some_0_tag_addr_is_garbage),
    .io_resp_bits_tag_addr_data(out_output_payload_Some_0_tag_addr_data),
    .io_resp_bits_tag_rows(out_output_payload_Some_0_tag_rows),
    .io_resp_bits_tag_cols(out_output_payload_Some_0_tag_cols),
    .io_resp_bits_data_0_0(out_output_payload_Some_0_data[0*20 +: 20]),
    .io_resp_bits_data_1_0(out_output_payload_Some_0_data[1*20 +: 20]),
    .io_resp_bits_data_2_0(out_output_payload_Some_0_data[2*20 +: 20]),
    .io_resp_bits_data_3_0(out_output_payload_Some_0_data[3*20 +: 20]),
    .io_resp_bits_data_4_0(out_output_payload_Some_0_data[4*20 +: 20]),
    .io_resp_bits_data_5_0(out_output_payload_Some_0_data[5*20 +: 20]),
    .io_resp_bits_data_6_0(out_output_payload_Some_0_data[6*20 +: 20]),
    .io_resp_bits_data_7_0(out_output_payload_Some_0_data[7*20 +: 20]),
    .io_resp_bits_data_8_0(out_output_payload_Some_0_data[8*20 +: 20]),
    .io_resp_bits_data_9_0(out_output_payload_Some_0_data[9*20 +: 20]),
    .io_resp_bits_data_10_0(out_output_payload_Some_0_data[10*20 +: 20]),
    .io_resp_bits_data_11_0(out_output_payload_Some_0_data[11*20 +: 20]),
    .io_resp_bits_data_12_0(out_output_payload_Some_0_data[12*20 +: 20]),
    .io_resp_bits_data_13_0(out_output_payload_Some_0_data[13*20 +: 20]),
    .io_resp_bits_data_14_0(out_output_payload_Some_0_data[14*20 +: 20]),
    .io_resp_bits_data_15_0(out_output_payload_Some_0_data[15*20 +: 20]),
    .io_resp_bits_total_rows(out_output_payload_Some_0_total_rows),
    .io_resp_bits_last(out_output_payload_Some_0_last),
    .io_tags_in_progress_0_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[0*1 +: 1]),
    .io_tags_in_progress_0_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[0*1 +: 1]),
    .io_tags_in_progress_0_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[0*1 +: 1]),
    .io_tags_in_progress_0_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[0*1 +: 1]),
    .io_tags_in_progress_0_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[0*1 +: 1]),
    .io_tags_in_progress_0_addr_data(in_input_0_3_resolver_inner_addr_data[0*14 +: 14]),
    .io_tags_in_progress_1_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[1*1 +: 1]),
    .io_tags_in_progress_1_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[1*1 +: 1]),
    .io_tags_in_progress_1_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[1*1 +: 1]),
    .io_tags_in_progress_1_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[1*1 +: 1]),
    .io_tags_in_progress_1_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[1*1 +: 1]),
    .io_tags_in_progress_1_addr_data(in_input_0_3_resolver_inner_addr_data[1*14 +: 14]),
    .io_tags_in_progress_2_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[2*1 +: 1]),
    .io_tags_in_progress_2_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[2*1 +: 1]),
    .io_tags_in_progress_2_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[2*1 +: 1]),
    .io_tags_in_progress_2_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[2*1 +: 1]),
    .io_tags_in_progress_2_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[2*1 +: 1]),
    .io_tags_in_progress_2_addr_data(in_input_0_3_resolver_inner_addr_data[2*14 +: 14]),
    .io_tags_in_progress_3_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[3*1 +: 1]),
    .io_tags_in_progress_3_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[3*1 +: 1]),
    .io_tags_in_progress_3_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[3*1 +: 1]),
    .io_tags_in_progress_3_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[3*1 +: 1]),
    .io_tags_in_progress_3_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[3*1 +: 1]),
    .io_tags_in_progress_3_addr_data(in_input_0_3_resolver_inner_addr_data[3*14 +: 14]),
    .io_tags_in_progress_4_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[4*1 +: 1]),
    .io_tags_in_progress_4_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[4*1 +: 1]),
    .io_tags_in_progress_4_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[4*1 +: 1]),
    .io_tags_in_progress_4_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[4*1 +: 1]),
    .io_tags_in_progress_4_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[4*1 +: 1]),
    .io_tags_in_progress_4_addr_data(in_input_0_3_resolver_inner_addr_data[4*14 +: 14]),
    .io_tags_in_progress_5_rob_id_valid(in_input_0_3_resolver_inner_rob_id_discriminant[5*1 +: 1]),
    .io_tags_in_progress_5_addr_is_acc_addr(in_input_0_3_resolver_inner_addr_is_acc_addr[5*1 +: 1]),
    .io_tags_in_progress_5_addr_accumulate(in_input_0_3_resolver_inner_addr_accumulate[5*1 +: 1]),
    .io_tags_in_progress_5_addr_read_full_acc_row(in_input_0_3_resolver_inner_addr_read_full_acc_row[5*1 +: 1]),
    .io_tags_in_progress_5_addr_garbage_bit(in_input_0_3_resolver_inner_addr_is_garbage[5*1 +: 1]),
    .io_tags_in_progress_5_addr_data(in_input_0_3_resolver_inner_addr_data[5*14 +: 14])
);

endmodule