module MeshWithDelaysBlackBoxAdapter(
    input           clock,
                    reset,
                    io_a_valid,
    input  [7:0]    io_a_bits_0_0,
                    io_a_bits_1_0,
                    io_a_bits_2_0,
                    io_a_bits_3_0,
                    io_a_bits_4_0,
                    io_a_bits_5_0,
                    io_a_bits_6_0,
                    io_a_bits_7_0,
                    io_a_bits_8_0,
                    io_a_bits_9_0,
                    io_a_bits_10_0,
                    io_a_bits_11_0,
                    io_a_bits_12_0,
                    io_a_bits_13_0,
                    io_a_bits_14_0,
                    io_a_bits_15_0,
    input           io_b_valid,
    input  [7:0]    io_b_bits_0_0,
                    io_b_bits_1_0,
                    io_b_bits_2_0,
                    io_b_bits_3_0,
                    io_b_bits_4_0,
                    io_b_bits_5_0,
                    io_b_bits_6_0,
                    io_b_bits_7_0,
                    io_b_bits_8_0,
                    io_b_bits_9_0,
                    io_b_bits_10_0,
                    io_b_bits_11_0,
                    io_b_bits_12_0,
                    io_b_bits_13_0,
                    io_b_bits_14_0,
                    io_b_bits_15_0,
    input           io_d_valid,
    input  [7:0]    io_d_bits_0_0,
                    io_d_bits_1_0,
                    io_d_bits_2_0,
                    io_d_bits_3_0,
                    io_d_bits_4_0,
                    io_d_bits_5_0,
                    io_d_bits_6_0,
                    io_d_bits_7_0,
                    io_d_bits_8_0,
                    io_d_bits_9_0,
                    io_d_bits_10_0,
                    io_d_bits_11_0,
                    io_d_bits_12_0,
                    io_d_bits_13_0,
                    io_d_bits_14_0,
                    io_d_bits_15_0,
    input           io_req_valid,
                    io_req_bits_tag_rob_id_valid,
    input  [5:0]    io_req_bits_tag_rob_id_bits,
    input           io_req_bits_tag_addr_is_acc_addr,
                    io_req_bits_tag_addr_accumulate,
                    io_req_bits_tag_addr_read_full_acc_row,
    input   [2:0]   io_req_bits_tag_addr_norm_cmd,              // DontCare
    input   [10:0]  io_req_bits_tag_addr_garbage,               // DontCare
                    io_req_bits_tag_addr_garbage_bit,
    input  [13:0]   io_req_bits_tag_addr_data,
    input  [4:0]    io_req_bits_tag_rows,
                    io_req_bits_tag_cols,
    input           io_req_bits_pe_control_dataflow,
                    io_req_bits_pe_control_propagate,
    input  [4:0]    io_req_bits_pe_control_shift,
    input           io_req_bits_a_transpose,
                    io_req_bits_bd_transpose,
    input  [4:0]    io_req_bits_total_rows,
    input  [1:0]    io_req_bits_flush,
    output          io_a_ready,
                    io_b_ready,
                    io_d_ready,
                    io_req_ready,
                    io_resp_valid,
                    io_resp_bits_tag_rob_id_valid,
    output [5:0]    io_resp_bits_tag_rob_id_bits,
    output          io_resp_bits_tag_addr_is_acc_addr,
                    io_resp_bits_tag_addr_accumulate,
                    io_resp_bits_tag_addr_read_full_acc_row,
    output [2:0]    io_resp_bits_tag_addr_norm_cmd,                     // DontCare
    output [10:0]   io_resp_bits_tag_addr_garbage,                      // DontCare
                    io_resp_bits_tag_addr_garbage_bit,
    output [13:0]   io_resp_bits_tag_addr_data,
    output [4:0]    io_resp_bits_tag_rows,
                    io_resp_bits_tag_cols,
    output [19:0]   io_resp_bits_data_0_0,
                    io_resp_bits_data_1_0,
                    io_resp_bits_data_2_0,
                    io_resp_bits_data_3_0,
                    io_resp_bits_data_4_0,
                    io_resp_bits_data_5_0,
                    io_resp_bits_data_6_0,
                    io_resp_bits_data_7_0,
                    io_resp_bits_data_8_0,
                    io_resp_bits_data_9_0,
                    io_resp_bits_data_10_0,
                    io_resp_bits_data_11_0,
                    io_resp_bits_data_12_0,
                    io_resp_bits_data_13_0,
                    io_resp_bits_data_14_0,
                    io_resp_bits_data_15_0,
    output [4:0]    io_resp_bits_total_rows,
    output          io_resp_bits_last,
                    io_tags_in_progress_0_rob_id_valid,
    output [5:0]    io_tags_in_progress_0_rob_id_bits,                    // DontCare
                    io_tags_in_progress_0_addr_is_acc_addr,
                    io_tags_in_progress_0_addr_accumulate,
                    io_tags_in_progress_0_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_0_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_0_addr_garbage,                   // DontCare
                    io_tags_in_progress_0_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_0_addr_data,
    output [4:0]    io_tags_in_progress_0_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_0_cols,                           // DontCare
    output          io_tags_in_progress_1_rob_id_valid,
    output [5:0]    io_tags_in_progress_1_rob_id_bits,                    // DontCare
                    io_tags_in_progress_1_addr_is_acc_addr,
                    io_tags_in_progress_1_addr_accumulate,
                    io_tags_in_progress_1_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_1_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_1_addr_garbage,                   // DontCare
                    io_tags_in_progress_1_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_1_addr_data,
    output [4:0]    io_tags_in_progress_1_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_1_cols,                           // DontCare
    output          io_tags_in_progress_2_rob_id_valid,
    output [5:0]    io_tags_in_progress_2_rob_id_bits,                    // DontCare
                    io_tags_in_progress_2_addr_is_acc_addr,
                    io_tags_in_progress_2_addr_accumulate,
                    io_tags_in_progress_2_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_2_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_2_addr_garbage,                   // DontCare
                    io_tags_in_progress_2_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_2_addr_data,
    output [4:0]    io_tags_in_progress_2_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_2_cols,                           // DontCare
    output          io_tags_in_progress_3_rob_id_valid,
    output [5:0]    io_tags_in_progress_3_rob_id_bits,                    // DontCare
                    io_tags_in_progress_3_addr_is_acc_addr,
                    io_tags_in_progress_3_addr_accumulate,
                    io_tags_in_progress_3_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_3_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_3_addr_garbage,                   // DontCare
                    io_tags_in_progress_3_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_3_addr_data,
    output [4:0]    io_tags_in_progress_3_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_3_cols,                           // DontCare
    output          io_tags_in_progress_4_rob_id_valid,
    output [5:0]    io_tags_in_progress_4_rob_id_bits,                    // DontCare
                    io_tags_in_progress_4_addr_is_acc_addr,
                    io_tags_in_progress_4_addr_accumulate,
                    io_tags_in_progress_4_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_4_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_4_addr_garbage,                   // DontCare
                    io_tags_in_progress_4_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_4_addr_data,
    output [4:0]    io_tags_in_progress_4_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_4_cols,                           // DontCare
    output          io_tags_in_progress_5_rob_id_valid,
    output [5:0]    io_tags_in_progress_5_rob_id_bits,                    // DontCare
                    io_tags_in_progress_5_addr_is_acc_addr,
                    io_tags_in_progress_5_addr_accumulate,
                    io_tags_in_progress_5_addr_read_full_acc_row,
    output [2:0]    io_tags_in_progress_5_addr_norm_cmd,                  // DontCare
    output [10:0]   io_tags_in_progress_5_addr_garbage,                   // DontCare
                    io_tags_in_progress_5_addr_garbage_bit,
    output [13:0]   io_tags_in_progress_5_addr_data,
    output [4:0]    io_tags_in_progress_5_rows,                           // DontCare
    output [4:0]    io_tags_in_progress_5_cols                            // DontCare
);
    wire [128-1:0] in_input_0_payload_Some_0_a_0;
    wire [128-1:0] in_input_1_payload_Some_0_b_0;
    wire [128-1:0] in_input_2_payload_Some_0_d_0;

    assign in_input_0_payload_Some_0_a_0[0*8 +: 8] = io_a_bits_0_0;
    assign in_input_0_payload_Some_0_a_0[1*8 +: 8] = io_a_bits_1_0;
    assign in_input_0_payload_Some_0_a_0[2*8 +: 8] = io_a_bits_2_0;
    assign in_input_0_payload_Some_0_a_0[3*8 +: 8] = io_a_bits_3_0;
    assign in_input_0_payload_Some_0_a_0[4*8 +: 8] = io_a_bits_4_0;
    assign in_input_0_payload_Some_0_a_0[5*8 +: 8] = io_a_bits_5_0;
    assign in_input_0_payload_Some_0_a_0[6*8 +: 8] = io_a_bits_6_0;
    assign in_input_0_payload_Some_0_a_0[7*8 +: 8] = io_a_bits_7_0;
    assign in_input_0_payload_Some_0_a_0[8*8 +: 8] = io_a_bits_8_0;
    assign in_input_0_payload_Some_0_a_0[9*8 +: 8] = io_a_bits_9_0;
    assign in_input_0_payload_Some_0_a_0[10*8 +: 8] = io_a_bits_10_0;
    assign in_input_0_payload_Some_0_a_0[11*8 +: 8] = io_a_bits_11_0;
    assign in_input_0_payload_Some_0_a_0[12*8 +: 8] = io_a_bits_12_0;
    assign in_input_0_payload_Some_0_a_0[13*8 +: 8] = io_a_bits_13_0;
    assign in_input_0_payload_Some_0_a_0[14*8 +: 8] = io_a_bits_14_0;
    assign in_input_0_payload_Some_0_a_0[15*8 +: 8] = io_a_bits_15_0;
    
    assign in_input_1_payload_Some_0_b_0[0*8 +: 8] = io_b_bits_0_0;
    assign in_input_1_payload_Some_0_b_0[1*8 +: 8] = io_b_bits_1_0;
    assign in_input_1_payload_Some_0_b_0[2*8 +: 8] = io_b_bits_2_0;
    assign in_input_1_payload_Some_0_b_0[3*8 +: 8] = io_b_bits_3_0;
    assign in_input_1_payload_Some_0_b_0[4*8 +: 8] = io_b_bits_4_0;
    assign in_input_1_payload_Some_0_b_0[5*8 +: 8] = io_b_bits_5_0;
    assign in_input_1_payload_Some_0_b_0[6*8 +: 8] = io_b_bits_6_0;
    assign in_input_1_payload_Some_0_b_0[7*8 +: 8] = io_b_bits_7_0;
    assign in_input_1_payload_Some_0_b_0[8*8 +: 8] = io_b_bits_8_0;
    assign in_input_1_payload_Some_0_b_0[9*8 +: 8] = io_b_bits_9_0;
    assign in_input_1_payload_Some_0_b_0[10*8 +: 8] = io_b_bits_10_0;
    assign in_input_1_payload_Some_0_b_0[11*8 +: 8] = io_b_bits_11_0;
    assign in_input_1_payload_Some_0_b_0[12*8 +: 8] = io_b_bits_12_0;
    assign in_input_1_payload_Some_0_b_0[13*8 +: 8] = io_b_bits_13_0;
    assign in_input_1_payload_Some_0_b_0[14*8 +: 8] = io_b_bits_14_0;
    assign in_input_1_payload_Some_0_b_0[15*8 +: 8] = io_b_bits_15_0;
    
    assign in_input_2_payload_Some_0_d_0[0*8 +: 8] = io_d_bits_0_0;
    assign in_input_2_payload_Some_0_d_0[1*8 +: 8] = io_d_bits_1_0;
    assign in_input_2_payload_Some_0_d_0[2*8 +: 8] = io_d_bits_2_0;
    assign in_input_2_payload_Some_0_d_0[3*8 +: 8] = io_d_bits_3_0;
    assign in_input_2_payload_Some_0_d_0[4*8 +: 8] = io_d_bits_4_0;
    assign in_input_2_payload_Some_0_d_0[5*8 +: 8] = io_d_bits_5_0;
    assign in_input_2_payload_Some_0_d_0[6*8 +: 8] = io_d_bits_6_0;
    assign in_input_2_payload_Some_0_d_0[7*8 +: 8] = io_d_bits_7_0;
    assign in_input_2_payload_Some_0_d_0[8*8 +: 8] = io_d_bits_8_0;
    assign in_input_2_payload_Some_0_d_0[9*8 +: 8] = io_d_bits_9_0;
    assign in_input_2_payload_Some_0_d_0[10*8 +: 8] = io_d_bits_10_0;
    assign in_input_2_payload_Some_0_d_0[11*8 +: 8] = io_d_bits_11_0;
    assign in_input_2_payload_Some_0_d_0[12*8 +: 8] = io_d_bits_12_0;
    assign in_input_2_payload_Some_0_d_0[13*8 +: 8] = io_d_bits_13_0;
    assign in_input_2_payload_Some_0_d_0[14*8 +: 8] = io_d_bits_14_0;
    assign in_input_2_payload_Some_0_d_0[15*8 +: 8] = io_d_bits_15_0;

    // Output wires.
    wire [320-1:0] out_output_payload_Some_0_data;

    // Resolver.
    wire [6-1:0] in_input_3_resolver_inner_rob_id_discriminant;
    wire [6-1:0] in_input_3_resolver_inner_addr_is_acc_addr;
    wire [6-1:0] in_input_3_resolver_inner_addr_accumulate;
    wire [6-1:0] in_input_3_resolver_inner_addr_read_full_acc_row;
    wire [6-1:0] in_input_3_resolver_inner_addr_is_garbage;
    wire [84-1:0] in_input_3_resolver_inner_addr_data;

    // DontCare resovler.
    wire [36-1:0] in_input_3_resolver_inner_rob_id_Some_0;
    wire [18-1:0] in_input_3_resolver_inner_addr_norm_cmd;
    wire [66-1:0] in_input_3_resolver_inner_addr_garbage;
    wire [30-1:0] in_input_3_resolver_inner_rows;
    wire [30-1:0] in_input_3_resolver_inner_cols;

    

    mwd_top mwd_inst(
        .clk(clock),
        .rst(reset),

        .in_input_0_payload_discriminant(io_a_valid),
        .in_input_0_payload_Some_0(in_input_0_payload_Some_0_a_0),
        .in_input_1_payload_discriminant(io_b_valid),
        .in_input_1_payload_Some_0(in_input_1_payload_Some_0_b_0),
        .in_input_2_payload_discriminant(io_d_valid),
        .in_input_2_payload_Some_0(in_input_2_payload_Some_0_d_0),
        .in_input_3_payload_discriminant(io_req_valid),
        .in_input_3_payload_Some_0_tag_rob_id_discriminant(io_req_bits_tag_rob_id_valid),
        .in_input_3_payload_Some_0_tag_rob_id_Some_0(io_req_bits_tag_rob_id_bits),
        .in_input_3_payload_Some_0_tag_addr_is_acc_addr(io_req_bits_tag_addr_is_acc_addr),
        .in_input_3_payload_Some_0_tag_addr_accumulate(io_req_bits_tag_addr_accumulate),
        .in_input_3_payload_Some_0_tag_addr_read_full_acc_row(io_req_bits_tag_addr_read_full_acc_row),
        .in_input_3_payload_Some_0_tag_addr_is_garbage(io_req_bits_tag_addr_garbage_bit),
        .in_input_3_payload_Some_0_tag_addr_data(io_req_bits_tag_addr_data),
        .in_input_3_payload_Some_0_tag_rows(io_req_bits_tag_rows),
        .in_input_3_payload_Some_0_tag_cols(io_req_bits_tag_cols),
        .in_input_3_payload_Some_0_pe_control_dataflow_discriminant(io_req_bits_pe_control_dataflow),
        .in_input_3_payload_Some_0_pe_control_propagate_discriminant(io_req_bits_pe_control_propagate),
        .in_input_3_payload_Some_0_pe_control_shift(io_req_bits_pe_control_shift),
        .in_input_3_payload_Some_0_transpose_a(io_req_bits_a_transpose),
        .in_input_3_payload_Some_0_transpose_bd(io_req_bits_bd_transpose),
        .in_input_3_payload_Some_0_total_rows(io_req_bits_total_rows),
        .in_input_3_payload_Some_0_flush(io_req_bits_flush),
        .in_input_3_payload_Some_0_tag_addr_norm_cmd(io_req_bits_tag_addr_norm_cmd),  // DontCare
        .in_input_3_payload_Some_0_tag_addr_garbage(io_req_bits_tag_addr_garbage),    // DontCare

        .in_input_0_resolver_ready(io_a_ready),
        .in_input_1_resolver_ready(io_b_ready),
        .in_input_2_resolver_ready(io_d_ready),
        .in_input_3_resolver_ready(io_req_ready),
        .in_input_3_resolver_inner_rob_id_discriminant(in_input_3_resolver_inner_rob_id_discriminant),
        .in_input_3_resolver_inner_rob_id_Some_0(in_input_3_resolver_inner_rob_id_Some_0), // Not used.
        .in_input_3_resolver_inner_addr_is_acc_addr(in_input_3_resolver_inner_addr_is_acc_addr),
        .in_input_3_resolver_inner_addr_accumulate(in_input_3_resolver_inner_addr_accumulate),
        .in_input_3_resolver_inner_addr_read_full_acc_row(in_input_3_resolver_inner_addr_read_full_acc_row),
        .in_input_3_resolver_inner_addr_norm_cmd(in_input_3_resolver_inner_addr_norm_cmd), // Not used.
        .in_input_3_resolver_inner_addr_garbage(in_input_3_resolver_inner_addr_garbage), // Not used.
        .in_input_3_resolver_inner_addr_is_garbage(in_input_3_resolver_inner_addr_is_garbage), 
        .in_input_3_resolver_inner_addr_data(in_input_3_resolver_inner_addr_data),
        .in_input_3_resolver_inner_rows(in_input_3_resolver_inner_rows), // Not used.
        .in_input_3_resolver_inner_cols(in_input_3_resolver_inner_cols), // Not used.

        .out_output_payload_discriminant(io_resp_valid),
        .out_output_payload_Some_0_tag_rob_id_discriminant(io_resp_bits_tag_rob_id_valid),
        .out_output_payload_Some_0_tag_rob_id_Some_0(io_resp_bits_tag_rob_id_bits),
        .out_output_payload_Some_0_tag_addr_is_acc_addr(io_resp_bits_tag_addr_is_acc_addr),
        .out_output_payload_Some_0_tag_addr_accumulate(io_resp_bits_tag_addr_accumulate),
        .out_output_payload_Some_0_tag_addr_read_full_acc_row(io_resp_bits_tag_addr_read_full_acc_row),
        .out_output_payload_Some_0_tag_addr_is_garbage(io_resp_bits_tag_addr_garbage_bit),
        .out_output_payload_Some_0_tag_addr_data(io_resp_bits_tag_addr_data),
        .out_output_payload_Some_0_tag_rows(io_resp_bits_tag_rows),
        .out_output_payload_Some_0_tag_cols(io_resp_bits_tag_cols),
        .out_output_payload_Some_0_data(out_output_payload_Some_0_data),
        .out_output_payload_Some_0_total_rows(io_resp_bits_total_rows),
        .out_output_payload_Some_0_last(io_resp_bits_last),

        .out_output_payload_Some_0_tag_addr_norm_cmd(io_resp_bits_tag_addr_norm_cmd), // Not used.
        .out_output_payload_Some_0_tag_addr_garbage(io_resp_bits_tag_addr_garbage) // Not used.
    );
    
    assign io_resp_bits_data_0_0 = out_output_payload_Some_0_data[0*20 +: 20];
    assign io_resp_bits_data_1_0 = out_output_payload_Some_0_data[1*20 +: 20];
    assign io_resp_bits_data_2_0 = out_output_payload_Some_0_data[2*20 +: 20];
    assign io_resp_bits_data_3_0 = out_output_payload_Some_0_data[3*20 +: 20];
    assign io_resp_bits_data_4_0 = out_output_payload_Some_0_data[4*20 +: 20];
    assign io_resp_bits_data_5_0 = out_output_payload_Some_0_data[5*20 +: 20];
    assign io_resp_bits_data_6_0 = out_output_payload_Some_0_data[6*20 +: 20];
    assign io_resp_bits_data_7_0 = out_output_payload_Some_0_data[7*20 +: 20];
    assign io_resp_bits_data_8_0 = out_output_payload_Some_0_data[8*20 +: 20];
    assign io_resp_bits_data_9_0 = out_output_payload_Some_0_data[9*20 +: 20];
    assign io_resp_bits_data_10_0 = out_output_payload_Some_0_data[10*20 +: 20];
    assign io_resp_bits_data_11_0 = out_output_payload_Some_0_data[11*20 +: 20];
    assign io_resp_bits_data_12_0 = out_output_payload_Some_0_data[12*20 +: 20];
    assign io_resp_bits_data_13_0 = out_output_payload_Some_0_data[13*20 +: 20];
    assign io_resp_bits_data_14_0 = out_output_payload_Some_0_data[14*20 +: 20];
    assign io_resp_bits_data_15_0 = out_output_payload_Some_0_data[15*20 +: 20];

    assign io_tags_in_progress_0_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[0];
    assign io_tags_in_progress_1_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[1];
    assign io_tags_in_progress_2_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[2];
    assign io_tags_in_progress_3_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[3];
    assign io_tags_in_progress_4_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[4];
    assign io_tags_in_progress_5_rob_id_valid = in_input_3_resolver_inner_rob_id_discriminant[5];

    assign io_tags_in_progress_0_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[0];
    assign io_tags_in_progress_1_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[1];
    assign io_tags_in_progress_2_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[2];
    assign io_tags_in_progress_3_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[3];
    assign io_tags_in_progress_4_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[4];
    assign io_tags_in_progress_5_addr_is_acc_addr = in_input_3_resolver_inner_addr_is_acc_addr[5];

    assign io_tags_in_progress_0_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[0];
    assign io_tags_in_progress_1_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[1];
    assign io_tags_in_progress_2_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[2];
    assign io_tags_in_progress_3_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[3];
    assign io_tags_in_progress_4_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[4];
    assign io_tags_in_progress_5_addr_accumulate = in_input_3_resolver_inner_addr_accumulate[5];

    assign io_tags_in_progress_0_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[0];
    assign io_tags_in_progress_1_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[1];
    assign io_tags_in_progress_2_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[2];
    assign io_tags_in_progress_3_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[3];
    assign io_tags_in_progress_4_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[4];
    assign io_tags_in_progress_5_addr_read_full_acc_row = in_input_3_resolver_inner_addr_read_full_acc_row[5];

    assign io_tags_in_progress_0_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[0];
    assign io_tags_in_progress_1_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[1];
    assign io_tags_in_progress_2_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[2];
    assign io_tags_in_progress_3_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[3];
    assign io_tags_in_progress_4_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[4];
    assign io_tags_in_progress_5_addr_garbage_bit = in_input_3_resolver_inner_addr_is_garbage[5];

    assign io_tags_in_progress_0_addr_data = in_input_3_resolver_inner_addr_data[0*14 +: 14];
    assign io_tags_in_progress_1_addr_data = in_input_3_resolver_inner_addr_data[1*14 +: 14];
    assign io_tags_in_progress_2_addr_data = in_input_3_resolver_inner_addr_data[2*14 +: 14];
    assign io_tags_in_progress_3_addr_data = in_input_3_resolver_inner_addr_data[3*14 +: 14];
    assign io_tags_in_progress_4_addr_data = in_input_3_resolver_inner_addr_data[4*14 +: 14];
    assign io_tags_in_progress_5_addr_data = in_input_3_resolver_inner_addr_data[5*14 +: 14];

    // DontCare

endmodule
    
                                 